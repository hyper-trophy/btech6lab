*U19Ec046 Resistively Loaded NMOS Inverter DC Analysis

.model mynmos nmos Vto=0.8 kp=20u

M1 out in 0 0 mynmos w=2u l=1u
Rl 1 out 200k
Vdd 1 0 5
Vin in 0 pulse (0 5 1ns 1ns 1ns 20ns 40ns)

.tran 1ns 50ns

.control
run
plot V(in) V(out)
.endc
.end