* U19EC046 Lab 2
.model mybjt npn (bf=20)
Q1 2 1 0 mybjt
Rc 2 3 1k
Rb 4 1 10k
Vcc 3 0 5
Vin 4 0 0

.dc Vin 0 5 0.05
.control
run
plot V(2) V(4)
.endc
.end


