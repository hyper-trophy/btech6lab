*CMOS Inverter

.model mynmos nmos Vto=0.8 Kp=50
.model mypmos pmos Vto=-1 Kp=20

Mn1 n_mn1_drain n_mn1_gate 0 0 mynmos w=1u l=1u
Mn2 n_mn1_drain n_mn2_gate 0 0 mynmos w=1u l=1u
Mp1 n_mp1_drain n_mn1_gate n_mp1_source n_mp1_source mypmos w=1.51u l=1u
Mp2 n_mn1_drain n_mn2_gate n_mp1_drain n_mp1_source mypmos w=1.51u l=1u

Mn3 n_mn2_gate n_mn3_gate 0 0 mynmos w=1u l=1u
Mn4 n_mn2_gate n_mn1_drain 0 0 mynmos w=1u l=1u
Mp3 n_mp3_drain n_mn3_gate n_mp1_source n_mp1_source mypmos w=1.51u l=1u
Mp4 n_mn2_gate n_mn1_drain n_mp3_drain n_mp1_source mypmos w=1.51u l=1u

Vdd n_mp1_source 0 5
* Vin1 n_mn1_gate 0 pulse(0 3 1ms 0 0 1ms 2ms)
* Vin2 n_mn3_gate 0 pulse(0 3 1ms 0 0 1ms 4ms)

Vin1 n_mn1_gate 0 5
Vin2 n_mn3_gate 0 5

.tran 1us 10ms

.control
run
* plot v(Va)
plot v(n_mn1_gate)
plot v(n_mn3_gate)
plot v(n_mn1_drain)
plot v(n_mn2_gate)
.endc
.end

* (5, 5, race, race), (0, 5, 5, 0), (5, 0, 0, 5), (0, 0, 2, 2)
*BICMOS transient char*

* .model q1 npn bf=50
* .model mynmos nmos Vto=0.8 Kp=50
* .model mypmos pmos Vto=-1 Kp=20

* .subckt BI in vdd_node out1 out2 src  
* M1 out1 in src src mynmos w=1u l=1u
* M2 out2 in vdd_node vdd_node mypmos w=1.51u l=1u
* .ends BI

* q11 vdd_node out2 out1 q1
* q12 out1 src 0 q1
* xd1 in1 vdd_node out1 out2 src BI
* Vdd vdd_node 0 5

* Vin in1 0 pulse(0 5 1ns 1ns 1ns 20us 40us)

* .tran 1ns 80us
* .control
* run
* plot v(in1) v(out1)
* .endc
* .end
