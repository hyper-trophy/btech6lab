* modified dtl propogation delay
.model mybjt npn bf=20
.model mydiode d

.subckt modifiedDTL in1 in2 vccNode gnd out
    rc vccNode out 2k
    q2 out q2base gnd mybjt
    r3 q2base gnd 5k
    dd q1emmiter q2base mydiode
    q1 q1collector q1base q1emmiter mybjt
    r2 q1collector q1base 2k
    r1 q1collector vccNode 1.75k
    da q1base in1 mydiode
    db q1base in2 mydiode
.ends dtlckt

*supply
vcc vccNode 0 5
* va in 0 pulse(0 5 0ps 10ps 10ps 200ps 1000ps)
va in 0 pulse(0 5 0ps 1ps 1ps 20us 40us)

Xd in in vccNode 0 out1 modifiedDTL
c_load out1 0 1p

.tran 20ns 80us

.control
run
plot v(in) v(out1)
.endc
.end