# CMOS
.model mynmos NMOS (Vt0=0.8, Kp=50u)
.model mypmos PMOS (Vt0=-1, Kp=20u)

.subckt cmosinverter in vdd_node out gnd
    MN out in gnd gnd mynmos w=1um l=50um
    MP vdd_node in out vdd_node mypmos w=2.5um l=50um
.ends cmosinverter

.subckt cmosinverter2 in vdd_node out gnd
    MN out in gnd gnd mynmos w=1um l=50um
    MP vdd_node in out vdd_node mypmos w=10um l=50um
.ends cmosinverter2

.subckt cmosinverter3 in vdd_node out gnd
    MN out in gnd gnd mynmos w=4um l=50um
    MP vdd_node in out vdd_node mypmos w=2.5um l=50um
.ends cmosinverter3


Vdd vdd_node 0 5
Vin input 0 5

Xd input vdd_node kr_0_25 0 cmosinverter
Xd2 input vdd_node kr_1 0 cmosinverter2
Xd3 input vdd_node kr_4 0 cmosinverter3

.dc Vin 0 5 0.005 

.control
run
plot v(input) v(kr_0_25) v(kr_1) v(kr_4)
.endc
.end
